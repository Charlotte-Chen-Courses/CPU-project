/////////////////////////////////////////////////////////////////////////
//                                                                     //
//   Modulename :  sys_defs.svh                                        //
//                                                                     //
//  Description :  This file has the macro-defines for macros used in  //
//                 the pipeline design.                                //
//                                                                     //
/////////////////////////////////////////////////////////////////////////

`ifndef __SYS_DEFS_SVH__
`define __SYS_DEFS_SVH__

// all files should `include "sys_defs.svh" to at least define the timescale
`timescale 1ns / 100ps

///////////////////////////////
// ---- Basic Constants ---- //
///////////////////////////////

// NOTE: the global CLOCK_PERIOD is defined in the Makefile

// useful boolean single-bit definitions
`define FALSE 1'h0
`define TRUE 1'h1

// data length
`define XLEN 32

// ROB number of entries
`define ROB_NUM_ENTRY 8

// RS number of entries
`define RS_NUM_ENTRY 5

// Map Table number of entries
`define MP_NUM_ENTRY 4

// CDB number of entries
`define CDB 2

// the zero register
// In RISC-V, any read of this register returns zero and any writes are thrown away
`define ZERO_REG 5'd0

// Basic NOP instruction. Allows pipline registers to clearly be reset with
// an instruction that does nothing instead of Zero which is really an ADDI x0, x0, 0
`define NOP 32'h00000013

//////////////////////////////////
// ---- Memory Definitions ---- //
//////////////////////////////////

// this will change for project 4
// the project 3 processor has a massive boost in performance just from having no mem latency
// see if you can beat it's CPI in project 4 even with a 100ns latency!
`define MEM_LATENCY_IN_CYCLES 0

`define NUM_MEM_TAGS 15

`define MEM_SIZE_IN_BYTES (64*1024)
`define MEM_64BIT_LINES (`MEM_SIZE_IN_BYTES/8)

typedef union packed {
  logic [7:0][7:0]  byte_level;
  logic [3:0][15:0] half_level;
  logic [1:0][31:0] word_level;
} EXAMPLE_CACHE_BLOCK;

typedef enum logic [1:0] {
  BYTE   = 2'h0,
  HALF   = 2'h1,
  WORD   = 2'h2,
  DOUBLE = 2'h3
} MEM_SIZE;

// Memory bus commands
typedef enum logic [1:0] {
  BUS_NONE  = 2'h0,
  BUS_LOAD  = 2'h1,
  BUS_STORE = 2'h2
} BUS_COMMAND;

///////////////////////////////
// ---- Exception Codes ---- //
///////////////////////////////

/**
 * Exception codes for when something goes wrong in the processor.
 * Note that we use HALTED_ON_WFI to signify the end of computation.
 * It's original meaning is to 'Wait For an Interrupt', but we generally
 * ignore interrupts in 470
 *
 * This mostly follows the RISC-V Privileged spec
 * except a few add-ons for our infrastructure
 * The majority of them won't be used, but it's good to know what they are
 */

typedef enum logic [3:0] {
  INST_ADDR_MISALIGN  = 4'h0,
  INST_ACCESS_FAULT   = 4'h1,
  ILLEGAL_INST        = 4'h2,
  BREAKPOINT          = 4'h3,
  LOAD_ADDR_MISALIGN  = 4'h4,
  LOAD_ACCESS_FAULT   = 4'h5,
  STORE_ADDR_MISALIGN = 4'h6,
  STORE_ACCESS_FAULT  = 4'h7,
  ECALL_U_MODE        = 4'h8,
  ECALL_S_MODE        = 4'h9,
  NO_ERROR            = 4'ha,  // a reserved code that we use to signal no errors
  ECALL_M_MODE        = 4'hb,
  INST_PAGE_FAULT     = 4'hc,
  LOAD_PAGE_FAULT     = 4'hd,
  HALTED_ON_WFI       = 4'he,  // 'Wait For Interrupt'. In 470, signifies the end of computation
  STORE_PAGE_FAULT    = 4'hf
} EXCEPTION_CODE;

////////////////////////////////////////
// ---- Datapath Control Signals ---- //
////////////////////////////////////////

// ALU opA input mux selects
typedef enum logic [1:0] {
  OPA_IS_RS1  = 2'h0,
  OPA_IS_NPC  = 2'h1,
  OPA_IS_PC   = 2'h2,
  OPA_IS_ZERO = 2'h3
} ALU_OPA_SELECT;

// ALU opB input mux selects
typedef enum logic [3:0] {
  OPB_IS_RS2   = 4'h0,
  OPB_IS_I_IMM = 4'h1,
  OPB_IS_S_IMM = 4'h2,
  OPB_IS_B_IMM = 4'h3,
  OPB_IS_U_IMM = 4'h4,
  OPB_IS_J_IMM = 4'h5
} ALU_OPB_SELECT;

// ALU function code input
// probably want to leave these alone
typedef enum logic [4:0] {
  ALU_ADD    = 5'h00,
  ALU_SUB    = 5'h01,
  ALU_SLT    = 5'h02,
  ALU_SLTU   = 5'h03,
  ALU_AND    = 5'h04,
  ALU_OR     = 5'h05,
  ALU_XOR    = 5'h06,
  ALU_SLL    = 5'h07,
  ALU_SRL    = 5'h08,
  ALU_SRA    = 5'h09,
  ALU_MUL    = 5'h0a,
  ALU_MULH   = 5'h0b,
  ALU_MULHSU = 5'h0c,
  ALU_MULHU  = 5'h0d,
  ALU_DIV    = 5'h0e,
  ALU_DIVU   = 5'h0f,
  ALU_REM    = 5'h10,
  ALU_REMU   = 5'h11
} FU_FUNC;

// Function Unit Marks
typedef enum logic [3:0] {
  ALU = 4'h0,
  LD  = 4'h1,
  ST  = 4'h2,
  FP1 = 4'h3,
  FP2 = 4'h4
} FUM;

// tag in map table
typedef enum logic [1:0] {
  REG_READY = 2'h0,  // value is ready in regfile
  NO_READY  = 2'h1,  // value is not ready
  ROB_READY = 4'h2   // value is ready in the ROB
  // we may need more bit
} TAG;

///////////////////////////////////
// ---- Instruction Typedef ---- //
///////////////////////////////////

typedef enum logic [2:0] {
  R = 3'h0,
  I = 3'h1,
  S = 3'h2,
  B = 3'h3,
  U = 3'h4,
  J = 3'h5
} INST_TYPE;

// from the RISC-V ISA spec
typedef union packed {
  logic [31:0] inst;
  INST_TYPE inst_type;
  struct packed {
    logic [6:0] funct7;
    logic [4:0] rs2;  // source register 2
    logic [4:0] rs1;  // source register 1
    logic [2:0] funct3;
    logic [4:0] rd;  // destination register
    logic [6:0] opcode;
  } r;  // register-to-register instructions
  struct packed {
    logic [11:0] imm;  // immediate value for calculating address
    logic [4:0] rs1;  // source register 1 (used as address base)
    logic [2:0] funct3;
    logic [4:0] rd;  // destination register
    logic [6:0] opcode;
  } i;  // immediate or load instructions
  struct packed {
    logic [6:0] off;  // offset[11:5] for calculating address
    logic [4:0] rs2;  // source register 2
    logic [4:0] rs1;  // source register 1 (used as address base)
    logic [2:0] funct3;
    logic [4:0] set;  // offset[4:0] for calculating address
    logic [6:0] opcode;
  } s;  // store instructions
  struct packed {
    logic       of;      // offset[12]
    logic [5:0] s;       // offset[10:5]
    logic [4:0] rs2;     // source register 2
    logic [4:0] rs1;     // source register 1
    logic [2:0] funct3;
    logic [3:0] et;      // offset[4:1]
    logic       f;       // offset[11]
    logic [6:0] opcode;
  } b;  // branch instructions
  struct packed {
    logic [19:0] imm;  // immediate value
    logic [4:0] rd;  // destination register
    logic [6:0] opcode;
  } u;  // upper-immediate instructions
  struct packed {
    logic       of;      // offset[20]
    logic [9:0] et;      // offset[10:1]
    logic       s;       // offset[11]
    logic [7:0] f;       // offset[19:12]
    logic [4:0] rd;      // destination register
    logic [6:0] opcode;
  } j;  // jump instructions

  // extensions for other instruction types
`ifdef ATOMIC_EXT
  struct packed {
    logic [4:0] funct5;
    logic       aq;
    logic       rl;
    logic [4:0] rs2;
    logic [4:0] rs1;
    logic [2:0] funct3;
    logic [4:0] rd;
    logic [6:0] opcode;
  } a;  // atomic instructions
`endif
`ifdef SYSTEM_EXT
  struct packed {
    logic [11:0] csr;
    logic [4:0]  rs1;
    logic [2:0]  funct3;
    logic [4:0]  rd;
    logic [6:0]  opcode;
  } sys;  // system call instructions
`endif

} INST;  // instruction typedef, this should cover all types of instructions


////////////////////////////////
// ---- Datapath Packets ---- //
////////////////////////////////

/**
 * Packets are used to move many variables between modules with
 * just one datatype, but can be cumbersome in some circumstances.
 *
 * Define new ones in project 4 at your own discretion
 */

/**
 * IF_DIS Packet:
 * Data exchanged from the IF to the Dispatch stage
 */
typedef struct packed {
  INST              inst;
  logic [`XLEN-1:0] PC;
  logic [`XLEN-1:0] NPC;    // PC + 4
  logic             valid;
} IF_DIS_PACKET;

/**
 * DIS_RM Packet:
 * Data exchanged from the Dispatch to the Rename stage
 */
typedef struct packed {
  INST              inst;
  logic [`XLEN-1:0] PC;
  logic [`XLEN-1:0] NPC;   // PC + 4

  logic [`XLEN-1:0] rs1_value;  // reg A value
  logic [`XLEN-1:0] rs2_value;  // reg B value

  ALU_OPA_SELECT opa_select;  // ALU opa mux select (ALU_OPA_xxx *)
  ALU_OPB_SELECT opb_select;  // ALU opb mux select (ALU_OPB_xxx *)

  logic [4:0] dest_reg_idx;  // destination (writeback) register index
  FU_FUNC fu_func;  // FU function select (ALU_xxx *)
  FUM fu_mark;  // FU function mark for RS
  logic rd_mem;  // Does inst read memory?
  logic wr_mem;  // Does inst write memory?
  logic cond_branch;  // Is inst a conditional branch?
  logic uncond_branch;  // Is inst an unconditional branch?
  logic pred_branch;  // Is inst an branch needs prediction
  logic halt;  // Is this a halt?
  logic illegal;  // Is this instruction illegal?
  logic csr_op;  // Is this a CSR operation? (we only used this as a cheap way to get return code)

  logic valid;
} DIS_RM_PACKET;



/**
 * RM_RSB Packet:
 * Data exchanged from the Dispatch to the Rename stage
 */
typedef struct packed {
  INST              inst;
  logic [`XLEN-1:0] PC;
  logic [`XLEN-1:0] NPC;   // PC + 4

  logic [`XLEN-1:0] rs1_value;  // reg A value
  logic [`XLEN-1:0] rs2_value;  // reg B value

  ALU_OPA_SELECT opa_select;  // ALU opa mux select (ALU_OPA_xxx *)
  ALU_OPB_SELECT opb_select;  // ALU opb mux select (ALU_OPB_xxx *)

  logic [4:0] dest_reg_idx;  // destination (writeback) register index
  FU_FUNC fu_func;  // FU function select (ALU_xxx *)
  FUM fu_mark;  // FU function mark for RS
  logic rd_mem;  // Does inst read memory?
  logic wr_mem;  // Does inst write memory?
  logic cond_branch;  // Is inst a conditional branch?
  logic uncond_branch;  // Is inst an unconditional branch?
  logic pred_branch;  // Is inst an branch needs prediction
  logic halt;  // Is this a halt?
  logic illegal;  // Is this instruction illegal?
  logic csr_op;  // Is this a CSR operation? (we only used this as a cheap way to get return code)

  logic valid;
} RM_RSB_PACKET;



/**
 * EX_MEM Packet:
 * Data exchanged from the EX to the MEM stage
 */
typedef struct packed {
  logic [`XLEN-1:0] alu_result;
  logic [`XLEN-1:0] NPC;

  logic             take_branch;   // Is this a taken branch?
  // Pass-through from decode stage
  logic [`XLEN-1:0] rs2_value;
  logic             rd_mem;
  logic             wr_mem;
  logic [4:0]       dest_reg_idx;
  logic             halt;
  logic             illegal;
  logic             csr_op;
  logic             rd_unsigned;   // Whether proc2Dmem_data is signed or unsigned
  MEM_SIZE          mem_size;
  logic             valid;
} EX_MEM_PACKET;

/**
 * MEM_WB Packet:
 * Data exchanged from the MEM to the WB stage
 *
 * Does not include data sent from the MEM stage to memory
 */
typedef struct packed {
  logic [`XLEN-1:0] result;
  logic [`XLEN-1:0] NPC;
  logic [4:0]       dest_reg_idx;  // writeback destination (ZERO_REG if no writeback)
  logic             take_branch;
  logic             halt;          // not used by wb stage
  logic             illegal;       // not used by wb stage
  logic             valid;
} MEM_WB_PACKET;

/**
 * No WB output packet as it would be more cumbersome than useful
 */

////////////////////////////////
// ------- OoO Entries ------ //
////////////////////////////////

/**
 * RS Entry:
 * Entries stored in Reservation Stations (RS)
 */
typedef struct packed {
  FUM               func_unit;          // functional unit mark for this entry
  logic             busy;               // If this functional unit is busy or not
  FU_FUNC           op_code;            // the operation of inst occupied this entry
  logic [4:0]       rob_target_index;   // index of this inst in ROB
  logic [4:0]       rob_source1_index;  // index of this first (left) reg of this inst in ROB
  logic [4:0]       rob_source2_index;  // index of this second (right) reg of this inst in ROB
  logic [`XLEN-1:0] source1_value;      // value in the first (left) reg of this inst
  logic             source1_ready;
  logic [`XLEN-1:0] source2_value;      // value in the second (right) reg of this inst
  logic             source2_ready;
  // we may need more entries
} RS_ENTRY;

/**
 * ROB Entry:
 * Entries stored in Reorder Buffer (ROB)
 */
typedef struct packed {
  logic [2:0]       ht;         // if this entry is head/tail
  logic [3:0]       index;      // entry index in ROB
  INST              inst;       // inst of this entry
  logic [4:0]       reg_index;  // target reg name of this inst
  logic [`XLEN-1:0] reg_value;  // value of the target reg
  // we may need more entries
} ROB_ENTRY;

/**
 * Map Table Entry:
 * Entries stored in Map Table (TB)
 */
typedef struct packed {
  logic [4:0] reg_index;  // reg name of this entry
  TAG         mp_tag;     // the status tag for this entry
  // we may need more entries
} TB_ENTRY;

/**
 * CDB Entry:
 * Entries for CDB broadcast
 */
typedef struct packed {
  logic [4:0]       rob_index;  // entry index in ROB
  logic [`XLEN-1:0] reg_value;  // value of the target reg in corresponding ROB entry
  // we may need more entries
} TB_ENTRY;


`endif  // __SYS_DEFS_SVH__
